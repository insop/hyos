--
-- package for tagged sorter: constant and others for 
--
-- Author: Insop Song
-- Begin Date  : 2007 05 01 
-- Ver   : 0.1
--
-- Revision History 
-- ---------------------------------------------------------------
-- Date         Author          Comments 
--
-- 
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

package tagged_pak is
    -- Design specific settings
    constant WIDTH_KEY  : integer := 32;
    constant WIDTH_DATA : integer := 32;
end tagged_pak;
